library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pc is
    port(
        rst: in std_logic;
        clk: in std_logic;
        wr_en: in std_logic;
        data_in: in unsigned(7 downto 0);
        data_out: out unsigned(7 downto 0):="00000000"
    );
end entity;

architecture a_pc of pc is
begin
    process(clk, rst)
    begin
        if rising_edge(clk) then
            if wr_en='1' and rst='0' then
                data_out<=data_in;
            end if;
        end if;
    end process;
end architecture;
